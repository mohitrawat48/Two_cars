/-------------------------------------------------------------------------
//      Two Cars Top Level   
//                                          
//      This is the top level,                                  
//      Set this file as top level before compilation                                   
//                                          
//      This module encompasses audio, keyboard and video subsystem                                    
//                                          
//                                          
//                                          
//                                          
//                                          
//-------------------------------------------------------------------------


module two_cars_top( input logic              CLOCK_50,
             input  logic      [3:0]  KEY,       
             output logic [6:0]  HEX0, HEX1,HEX2,HEX3,HEX4,HEX5,HEX6,HEX7,
				 output logic [2:0] LEDG,
             // VGA Interface 
             output logic [7:0]  VGA_R,        //VGA Red
                                 VGA_G,        //VGA Green
                                 VGA_B,        //VGA Blue
             output logic        VGA_CLK,      //VGA Clock
                                 VGA_SYNC_N,   //VGA Sync signal
                                 VGA_BLANK_N,  //VGA Blank signal
                                 VGA_VS,       //VGA virtical sync signal
                                 VGA_HS,       //VGA horizontal sync signal
											
             // CY7C67200 Interface
             inout  wire  [15:0] OTG_DATA,     //CY7C67200 Data bus 16 Bits
             output logic [1:0]  OTG_ADDR,     //CY7C67200 Address 2 Bits
             output logic        OTG_CS_N,     //CY7C67200 Chip Select
                                 OTG_RD_N,     //CY7C67200 Write
                                 OTG_WR_N,     //CY7C67200 Read
                                 OTG_RST_N,    //CY7C67200 Reset
             input               OTG_INT,      //CY7C67200 Interrupt
				 
             // SDRAM Interface for Nios II Software
             output logic [12:0] DRAM_ADDR,    //SDRAM Address 13 Bits
             inout  wire  [31:0] DRAM_DQ,      //SDRAM Data 32 Bits
             output logic [1:0]  DRAM_BA,      //SDRAM Bank Address 2 Bits
             output logic [3:0]  DRAM_DQM,     //SDRAM Data Mast 4 Bits
             output logic        DRAM_RAS_N,   //SDRAM Row Address Strobe
                                 DRAM_CAS_N,   //SDRAM Column Address Strobe
                                 DRAM_CKE,     //SDRAM Clock Enable
                                 DRAM_WE_N,    //SDRAM Write Enable
                                 DRAM_CS_N,    //SDRAM Chip Select
                                 DRAM_CLK,      //SDRAM Clock
             //SRAM Signals
				 output logic SRAM_CE_N, SRAM_UB_N, SRAM_LB_N, SRAM_OE_N, SRAM_WE_N,
             output logic [19:0] SRAM_ADDR,
             inout wire [15:0] SRAM_DQ,
				 
				 
				 //audio signals
				   //audio chip
				 input logic AUD_ADCDAT, AUD_DACLRCK, AUD_ADCLRCK, AUD_BCLK,
				 output logic AUD_DACDAT, AUD_XCK, I2C_SCLK, I2C_SDAT,
					//flash memory
				 output logic [22:0] FL_ADDR,
				 input logic [7:0] FL_DQ,
				 output logic FL_WE_N,FL_RST_N,FL_WP_N,FL_CE_N,FL_OE_N
				 );
						  
	 //We wanted to run Sram as fast as poosible
	 //It can be run at Maximum of 100Mhz
	 //Sram has seprate Clk
	 //this 100Mhz clock is generated by a PLL module in Qsys
	 logic sram_clk;
	 
	 // Reset_h  resets the audio
	 // Reset_h1 resets the game
    logic Reset_h,Reset_h1, Clk;
    logic [15:0] keycode;
    
    assign Clk = CLOCK_50;
    always_ff @ (posedge Clk) begin
        Reset_h <= ~(KEY[0]);        // The push buttons are active low
		  Reset_h1 <= ~(KEY[1]);
    end
    
	 
	 
    // Interface signals between NIOS II and EZ-OTG chip
    logic [1:0] hpi_addr;
    logic [15:0] hpi_data_in, hpi_data_out;
    logic hpi_r, hpi_w, hpi_cs, hpi_reset;
    
    // Interface between NIOS II and EZ-OTG chip
    hpi_io_intf hpi_io_inst(
                            .Clk(Clk),
                            .Reset(Reset_h1),
                            // signals connected to NIOS II
                            .from_sw_address(hpi_addr),
                            .from_sw_data_in(hpi_data_in),
                            .from_sw_data_out(hpi_data_out),
                            .from_sw_r(hpi_r),
                            .from_sw_w(hpi_w),
                            .from_sw_cs(hpi_cs),
                            .from_sw_reset(hpi_reset),
                            // signals connected to EZ-OTG chip
                            .OTG_DATA(OTG_DATA),    
                            .OTG_ADDR(OTG_ADDR),    
                            .OTG_RD_N(OTG_RD_N),    
                            .OTG_WR_N(OTG_WR_N),    
                            .OTG_CS_N(OTG_CS_N),
                            .OTG_RST_N(OTG_RST_N)
    );
     
     // You need to make sure that the port names here match the ports in Qsys-generated codes.
     lab8_soc my_lab8_soc(        //modified line orig: nios_system nios_system
                             .clk_clk(Clk),         
                             .reset_reset_n(1'b1),    // Never reset NIOS
                             .sdram_wire_addr(DRAM_ADDR), 
                             .sdram_wire_ba(DRAM_BA),   
                             .sdram_wire_cas_n(DRAM_CAS_N),
                             .sdram_wire_cke(DRAM_CKE),  
                             .sdram_wire_cs_n(DRAM_CS_N), 
                             .sdram_wire_dq(DRAM_DQ),   
                             .sdram_wire_dqm(DRAM_DQM),  
                             .sdram_wire_ras_n(DRAM_RAS_N),
                             .sdram_wire_we_n(DRAM_WE_N), 
                             .sdram_clk_clk(DRAM_CLK),
                             .keycode_export(keycode),  
                             .otg_hpi_address_export(hpi_addr),
                             .otg_hpi_data_in_port(hpi_data_in),
                             .otg_hpi_data_out_port(hpi_data_out),
                             .otg_hpi_cs_export(hpi_cs),
                             .otg_hpi_r_export(hpi_r),
                             .otg_hpi_w_export(hpi_w),
                             .otg_hpi_reset_export(hpi_reset),
									  .sram_clk_clk(sram_clk)
    );

	
 
    // PLL has been to to generate the 25MHZ VGA_CLK.
	 // VGA runs at 25 Mhz,
    vga_clk vga_clk_instance(.inclk0(Clk), .c0(VGA_CLK));
    
	 
	 //VGA signals for intermodule connection
	 logic [9:0] my_DrawX,my_DrawY;
	 logic my_VGA_VS;
	 assign VGA_VS = my_VGA_VS;
	 
	 //signals for intermodule connection 
	 logic [7:0] player1_key, player2_key;
	 
	 //VGA controller 
	 //generates VGA control signals
	 VGA_controller vga_controller_instance(.Clk(Clk), .Reset(Reset_h1), 
								.VGA_CLK(VGA_CLK),.VGA_HS(VGA_HS),.VGA_VS(my_VGA_VS), 
								.VGA_BLANK_N(VGA_BLANK_N),.VGA_SYNC_N(VGA_SYNC_N),
								.DrawX(my_DrawX), .DrawY(my_DrawY));
	 

	  //The purpose of this signal is to check 'Enter' Keypress
	  //User Presses Enter Key to exit Menu screen and start the game
	  logic [7:0] keys;
	  assign keys = keycode[7:0];
	 
	 //This module literaly contains the entire game mechanics
	 //Everthing except keyboard and audio is inside this module
	 VGA_manager my_VGA_manager( .*,.Clk(sram_clk), .Reset(Reset_h1),.frame_clk(my_VGA_VS),
										  .VGA_R(VGA_R),.VGA_G(VGA_G),.VGA_B(VGA_B),
								        .X_Cord(my_DrawX),.Y_Cord(my_DrawY),
										  .CE(SRAM_CE_N),.UB(SRAM_UB_N),
										  .LB(SRAM_LB_N),.OE(SRAM_OE_N),.WE(SRAM_WE_N),
										  .ADDR(SRAM_ADDR),.Data(SRAM_DQ),.keycode(keys) 
								        );
	 
	 
	 //This module takes two keypresses from NIOS at a time 
	 //and separates them into two groups player1_key and player2_key
	 mapkeys my_map_keys( .player1_key(player1_key), .player2_key(player2_key),
								 .two_keycodes(keycode) );
		
	 //fecthes data from flash memory and sends to audio chip
	 audio_monitor my_audio_machine(.*,.Reset(Reset_h));
	 
    // Display player1 and player2 keypresses on hex display
    HexDriver hex_inst_0 (player2_key[3:0], HEX0);
    HexDriver hex_inst_1 (player2_key[7:4], HEX1);
	 HexDriver hex_inst_2 (player1_key[3:0], HEX2);
	 HexDriver hex_inst_3 (player1_key[7:4], HEX3);
	 
	 //Displays keypresses from NIOS on hex display
    HexDriver hex_inst_4 (keycode[3:0], HEX4);
    HexDriver hex_inst_5 (keycode[7:4], HEX5);
	 HexDriver hex_inst_6 (keycode[11:8], HEX6);
	 HexDriver hex_inst_7 (keycode[15:12], HEX7);
 
 
endmodule
